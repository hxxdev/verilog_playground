`ifndef ALU_TB_PKG_SV
`define ALU_TB_PKG_SV

package alu_tb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "alu_transaction.sv"
  `include "alu_driver.sv"
  `include "alu_monitor.sv"
  `include "alu_scoreboard.sv"
  `include "alu_env.sv"
  `include "alu_test.sv"

endpackage

`endif
