module top ();

  counter u_counter (
      .i_clk(),
      .clk(),
      .en(en),
      .rst(rst),
      .count(count)
  );

  initial begin

  end

endmodule
