module top ();
    counter u_counter (
        .clk(),
        .en(),
        .rst(),
        .count(),
    );
endmodule
